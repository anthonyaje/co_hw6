//Subject:     CO project 2 - PC
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Luke
//----------------------------------------------
//Date:        2010/8/16
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module ProgramCounter(
    clk_i,
	rst_n,
	pc_in_i,
	pc_load_control,
	pc_out_o
	);
     
//I/O ports
input           clk_i;
input	        rst_n;
input 			pc_load_control;
input  [32-1:0] pc_in_i;
output [32-1:0] pc_out_o;
 
//Internal Signals
reg    [32-1:0] pc_out_o;
 
//Parameter

    
//Main function
always @(posedge clk_i) begin
    if(~rst_n)
	    pc_out_o <= 0;
	else if(pc_load_control)begin
		//do nothing
	end
	else
	    pc_out_o <= pc_in_i;
end

endmodule



                    
                    